module InstructionFetch(
			input );
   
endmodule
