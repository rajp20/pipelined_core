module InstructionFetch(
			input 		  clk,
			input      [15:0] PC,
			input      [15:0] TARGET, 
			input      [15:0] data_from_mem,
			output reg [15:0] NPC_IF,
			output reg [15:0] INST_IF);

   
endmodule
