module InstructionDecode(input             clk,
			 input      [15:0] NPC_IF,
			 input      [15:0] INST_IF,
			 output reg [15:0] NPC_ID,
			 output reg [15:0] REG1_ID
			 output reg [15:0] REG2_ID
			 output reg [4:0]  CTRL_ID);

endmodule
