module InstructionFetch(input 		  clk,
			input [15:0] 	  PC,
			input [15:0] 	  TARGET,
			input 		  TARGET_EN, 
			input [15:0] 	  from_mem_data,
			output reg [15:0] to_mem_addr,
			output reg [15:0] NPC_IF,
			output reg [15:0] INST_IF);

   
endmodule
